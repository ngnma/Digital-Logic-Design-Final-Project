module f1_tb ();
	reg a,a2,b,b2,c,c2,d,d2;
	wire out;
	f1 f1(out,a,a2,b,b2,c,c2,d,d2);
	initial begin
			$dumpfile("f1.vcd");
			$dumpvars(0,f1_tb);
			a=0;
			b=0;
			c=0;
			d=0;
			a2=1;
			b2=1;
			c2=1;
			d2=1;
			#20;
			a=1;
			a2=0;
			#20;
			b=1;
			b2=0;
			#20;
			a=0;
			a2=1;
			#20;
			c=1;
			c2=0;
			#20;
			a=1;
			a2=0;
			#20;
			b=0;
			b2=1;
			#20;
			a=0;
			a2=1;
			#20;
			d=1;
			d2=0;
			#20;
			a=1;
			a2=0;
			#20;
			b=1;
			b2=0;
			#20;
			a=0;
			a2=1;
			#20;
			c=0;
			c2=1;
			#20;
			a=1;
			a2=0;
			#20;
			b=0;
			b2=1;
			#20;
			a=0;
			a2=1;
			#20;
		end

endmodule